-- Listing 13.7
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity pong_graph is
   port(
      clk, reset: std_logic;
      btn: std_logic_vector(3 downto 0);
		shoot, d_clr: std_logic; --switch1
      pixel_x,pixel_y: in std_logic_vector(9 downto 0);
      gra_still, d_inc: in std_logic;
		--dig0: in std_logic_vector(3 downto 0);
      --graph_on, hit, miss: out std_logic;
		graph_on, miss: out std_logic;
      rgb: out std_logic_vector(2 downto 0);
		hiteI,hiteII,hiteIII: out std_logic;
		rst_enemy: in std_logic_vector(2 downto 0);
		arrows: in std_logic_vector(4 downto 0)
   );
end pong_graph;

architecture arch of pong_graph is
   signal pix_x, pix_y: unsigned(9 downto 0);
	signal btn_reg, btn_next: std_logic_vector(3 downto 0);
	signal arrow_reg, arrow_next: std_logic_vector(4 downto 0);
   constant MAX_X: integer:=640;
   constant MAX_Y: integer:=480;
	constant zero: integer:= 0;
	constant eight: integer:=8;
	
	signal shot_next,shot_reg: std_logic := '0';
	
	--constant CHESS_SQR: integer := 32;
   
	--constant WALL_X_L_L: integer:=0;
   --constant WALL_X_R_L: integer:=8;
	--constant WALL_X_L_R: integer:=630;
   --constant WALL_X_R_R: integer:=640;
	
	--constant WALL_Y_T_T: integer:=0;
	--constant WALL_Y_B_T: integer:=8;
	--constant WALL_Y_T_B: integer:=456-9; -- 480 - 
	--constant WALL_Y_B_B: integer:=480;
	
   signal player_y_t, player_y_b, player_x_r, player_x_l: unsigned(9 downto 0);
   --constant PLAYER_SIZE: integer:=32;
	--constant PLAYER_X_Size: integer:=32;
   signal player_y_reg, player_y_next: unsigned(9 downto 0);
	signal player_x_reg, player_x_next: unsigned(9 downto 0);
   constant PLAYER_V: integer:=2;
   --constant BALL_SIZE: integer:=8; -- 8
   signal ball_x_l, ball_x_r: unsigned(9 downto 0);
   signal ball_y_t, ball_y_b: unsigned(9 downto 0);
   signal ball_x_reg, ball_x_next: unsigned(9 downto 0);
   signal ball_y_reg, ball_y_next: unsigned(9 downto 0);
   signal ball_vx_reg, ball_vx_next: unsigned(9 downto 0);
   signal ball_vy_reg, ball_vy_next: unsigned(9 downto 0);
   constant BALL_V_P: unsigned(9 downto 0)
            :=to_unsigned(4,10);
   constant BALL_V_N: unsigned(9 downto 0)
            :=unsigned(to_signed(-4,10));
	--constant BALL_V_Z: unsigned(9 downto 0)
   --         :=unsigned(to_signed(0,10));
				
				
--ENEMY ----------------------------------------------------------				
	constant ENEMY_SIZE: integer:=32;
	--constant ENEMY_X_SIZE: integer:=32;
	constant ENEMY_V_P: unsigned(9 downto 0)
            :=to_unsigned(1,10);
   constant ENEMY_V_N: unsigned(9 downto 0)
            :=unsigned(to_signed(-1,10));
	constant ENEMY_V_Z: unsigned(9 downto 0)
            :=unsigned(to_signed(0,10));	
				
   signal enemy_x_l, enemy_x_r: unsigned(9 downto 0);
   signal enemy_y_t, enemy_y_b: unsigned(9 downto 0);
   signal enemy_x_reg, enemy_x_next: unsigned(9 downto 0);
   signal enemy_y_reg, enemy_y_next: unsigned(9 downto 0);
   signal enemy_vx_reg, enemy_vx_next: unsigned(9 downto 0);
   signal enemy_vy_reg, enemy_vy_next: unsigned(9 downto 0);
	
	signal enemyII_x_l, enemyII_x_r: unsigned(9 downto 0);
   signal enemyII_y_t, enemyII_y_b: unsigned(9 downto 0);
   signal enemyII_x_reg, enemyII_x_next: unsigned(9 downto 0);
   signal enemyII_y_reg, enemyII_y_next: unsigned(9 downto 0);
   signal enemyII_vx_reg, enemyII_vx_next: unsigned(9 downto 0);
   signal enemyII_vy_reg, enemyII_vy_next: unsigned(9 downto 0);
	
	signal enemyIII_x_l, enemyIII_x_r: unsigned(9 downto 0);
   signal enemyIII_y_t, enemyIII_y_b: unsigned(9 downto 0);
   signal enemyIII_x_reg, enemyIII_x_next: unsigned(9 downto 0);
   signal enemyIII_y_reg, enemyIII_y_next: unsigned(9 downto 0);
   signal enemyIII_vx_reg, enemyIII_vx_next: unsigned(9 downto 0);
   signal enemyIII_vy_reg, enemyIII_vy_next: unsigned(9 downto 0);
	
				
--BULLET-----------------------------------------------------------
   type rom_type is array (0 to 7) of
        std_logic_vector (7 downto 0);
   constant BALL_ROM: rom_type :=
   (
      "00000000", --   ****
      "00111100", --  ******
      "01111110", -- ********
      "11111111", -- ********
      "11111111", -- ********
      "01111110", -- ********
      "00111100", --  ******
      "00000000"  --   ****
   );
-------------------------------------------------------------------
	type rom_type_2 is array (0 to 31, 0 to 31) of std_logic_vector (2 downto 0);
	constant PLAYER_ROM: rom_type_2 :=
   (
       ("000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "001", "001", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "001", "001", "110", "110", "001", "001", "001", "110", "110", "110", "110", "001", "001", "001", "110", "110", "001", "001", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "001", "001", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "001", "001", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "001", "001", "110", "110", "110", "110", "000", "001", "110", "110", "110", "110", "001", "000", "110", "110", "110", "110", "001", "001", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "001", "001", "110", "110", "110", "110", "000", "001", "110", "110", "110", "110", "001", "000", "110", "110", "110", "110", "001", "001", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "001", "001", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "001", "001", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "001", "001", "000", "000", "000", "000", "011", "011", "011", "011", "011", "011", "011", "011", "000", "000", "000", "000", "001", "001", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "001", "110", "110", "110", "110", "011", "011", "011", "011", "011", "011", "011", "011", "110", "110", "110", "110", "001", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "011", "011", "011", "011", "011", "011", "011", "011", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "011", "011", "011", "011", "011", "011", "011", "011", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "010", "010", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "010", "010", "010", "010", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "001", "010", "101", "101", "010", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "110", "110", "010", "101", "101", "010", "110", "110", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "110", "110", "010", "010", "010", "010", "110", "110", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "110", "110", "110", "110", "110", "110", "110", "110", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "110", "110", "110", "110", "110", "110", "110", "110", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "100", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000")
   );
	
	constant PLAYER_ROM_SIDE: rom_type_2 :=
   (
       ("000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "001", "001", "001", "001", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "001", "001", "001", "001", "001", "110", "110", "001", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "001", "001", "001", "001", "001", "001", "001", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "101", "101", "101", "001", "001", "001", "001", "001", "001", "001", "001", "110", "110", "110", "110", "000", "001", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "001", "001", "001", "001", "110", "110", "110", "001", "001", "001", "110", "110", "110", "110", "110", "000", "001", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "001", "001", "001", "001", "110", "110", "110", "110", "110", "001", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "001", "001", "001", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "011", "011", "011", "011", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "001", "110", "110", "110", "110", "000", "110", "110", "110", "110", "110", "110", "110", "011", "011", "011", "011", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "000", "110", "110", "110", "110", "110", "110", "110", "011", "011", "011", "011", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "011", "011", "011", "011", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "010", "010", "010", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "010", "010", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "010", "000", "000"),
		 ("000", "000", "000", "011", "011", "000", "010", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "010", "010", "010", "010", "010", "000", "000"),
		 ("000", "000", "000", "011", "011", "011", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "010", "010", "010", "010", "010", "000", "000"),
		 ("000", "000", "000", "011", "011", "011", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "110", "110", "010", "010", "010", "010", "000", "000"),
		 ("000", "000", "000", "011", "011", "011", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "110", "110", "010", "010", "000", "000", "000", "000"),
		 ("000", "000", "000", "011", "011", "011", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "001", "001", "001", "001", "001", "110", "110", "110", "110", "000", "000", "000", "000"),
		 ("000", "000", "000", "011", "011", "011", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "001", "001", "001", "001", "110", "110", "110", "110", "000", "000", "000", "000"),
		 ("000", "000", "000", "011", "011", "011", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "001", "001", "100", "100", "100", "100", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "100", "100", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000")
   );
	
	constant PLAYER_ROM_BACK: rom_type_2 :=
   (
       ("000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "001", "001", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "001", "001", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "001", "001", "001", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "001", "001", "001", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "001", "001", "001", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "101", "001", "001", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "110", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "010", "010", "010", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "010", "010", "010", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "010", "010", "000", "000", "000", "000", "000", "000", "000", "000", "010", "010", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "010", "000", "000", "000", "000", "000", "011", "011", "011", "010", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "011", "000", "000", "011", "011", "011", "011", "011", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "011", "011", "011", "011", "011", "011", "011", "011", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "011", "011", "011", "011", "011", "011", "011", "011", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "011", "011", "011", "011", "011", "011", "011", "011", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "011", "011", "011", "011", "011", "011", "011", "011", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "011", "011", "011", "011", "011", "011", "011", "011", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "000", "100", "100", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000"),
		 ("000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000", "000")
   );
	type rom_type_3 is array (0 to 15,0 to 15) of
        std_logic_vector (2 downto 0);
	constant ENEMY_ROM_SIDE: rom_type_3 :=
	(
		("000","000", "000", "000", "001", "000", "000", "001", "000", "001", "001", "000", "000", "000", "000", "000"),
		("000","000", "000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000", "000"),
		("000","000", "000", "001", "001", "001", "001", "001", "001", "001", "001", "001", "001", "000", "000", "000"),
		("000","000", "000", "000", "001", "001", "110", "110", "001", "001", "110", "001", "000", "000", "000", "000"),
		("000","000", "000", "001", "001", "001", "110", "110", "110", "110", "110", "100", "000", "000", "000", "000"),
		("000","000", "000", "001", "001", "110", "110", "110", "110", "110", "010", "110", "000", "000", "000", "000"),
		("000","000", "000", "000", "001", "110", "110", "110", "110", "110", "110", "010", "000", "000", "000", "000"),
		("000","000", "000", "000", "000", "010", "100", "100", "100", "100", "100", "011", "100", "110", "000", "000"),
		("000","000", "000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000"),
		("000","000", "000", "000", "011", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "110"),
		("000","000", "000", "000", "011", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000"),
		("000","000", "000", "000", "011", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000"),
		("000","000", "000", "000", "100", "100", "100", "100", "100", "100", "100", "100", "000", "000", "000", "000"),
		("000","000", "000", "000", "000", "001", "100", "000", "000", "100", "100", "100", "100", "000", "000", "000"),
		("000","000", "000", "000", "000", "001", "001", "000", "000", "000", "001", "001", "000", "000", "000", "000"),
		("000","000", "000", "000", "000", "000", "001", "001", "000", "000", "001", "001", "001", "000", "000", "000")
	);
	
   
	signal rom_addr_player, rom_col_player: unsigned(5 downto 0);
	signal rom_bit_player,rom_next_player: std_logic_vector(2 downto 0);
	--signal rom_data_player: std_logic_vector(7 downto 0);
	
	signal rom_addr_enemy, rom_col_enemy: unsigned(3 downto 0);
	signal rom_bit_enemy, rom_next_enemy: std_logic_vector(2 downto 0);
	--signal rom_data_enemy: std_logic_vector(7 downto 0);
	
	signal rom_addr_enemyII, rom_col_enemyII: unsigned(3 downto 0);
	signal rom_bit_enemyII, rom_next_enemyII: std_logic_vector(2 downto 0);
	--signal rom_data_enemyII: std_logic_vector(7 downto 0);
	
	signal rom_addr_enemyIII, rom_col_enemyIII: unsigned(3 downto 0);
	signal rom_bit_enemyIII, rom_next_enemyIII: std_logic_vector(2 downto 0);
	--signal rom_data_enemyIII: std_logic_vector(7 downto 0);
	
	signal rom_addr, rom_col: unsigned(2 downto 0);
   signal rom_data: std_logic_vector(7 downto 0);
   signal rom_bit: std_logic;
   signal wall_on, rd_ball_on, player_on, enemy_on, enemyII_on, enemyIII_on: std_logic;

   signal wall_rgb, player_rgb, ball_rgb, enemy_rgb, enemyII_rgb, enemyIII_rgb:std_logic_vector(2 downto 0);
   signal refr_tick: std_logic;
	signal contador,contador_next: std_logic_vector(1 downto 0);

	
begin
	-----------------------------------------------------------
   -- REGISTERS
	-----------------------------------------------------------
   process (clk,reset)
   begin
      if reset='1' then
		
         player_y_reg <= (OTHERS=>'0');
			player_x_reg <= (OTHERS=>'0');
         
			ball_x_reg <= (OTHERS=>'0');
         ball_y_reg <= (OTHERS=>'0');
         ball_vx_reg <= ("0000000100");
         ball_vy_reg <= ("0000000100");
			
			enemy_x_reg <= (OTHERS=>'0');
         enemy_y_reg <= (OTHERS=>'0');
         enemy_vx_reg <= ("0000000100");
         enemy_vy_reg <= ("0000000100");
			
			enemyII_x_reg <= (OTHERS=>'0');
         enemyII_y_reg <= (OTHERS=>'0');
         enemyII_vx_reg <= ("0000000100");
         enemyII_vy_reg <= ("0000000100");
			
			enemyIII_x_reg <= (OTHERS=>'0');
			enemyIII_y_reg <= (OTHERS=>'0');
			enemyIII_vx_reg <= ("0000000100");
			enemyIII_vy_reg <= ("0000000100");
			
			shot_reg <= '0';
			rom_bit_player <= (OTHERS=>'0');
			btn_reg <= (others=>'0');
			arrow_reg <=(others =>'0');
			
			rom_bit_enemy <= (OTHERS => '0');
			rom_bit_enemyII <= (OTHERS => '0');
			rom_bit_enemyIII <= (OTHERS => '0');
			contador <= (OTHERS => '0');
      elsif (clk'event and clk='1') then
		
         player_y_reg <= player_y_next;
			player_x_reg <= player_x_next;
			
         ball_x_reg <= ball_x_next;
         ball_y_reg <= ball_y_next;
         ball_vx_reg <= ball_vx_next;
         ball_vy_reg <= ball_vy_next;
			
			enemy_x_reg <= enemy_x_next;
         enemy_y_reg <= enemy_y_next;
         enemy_vx_reg <= enemy_vx_next;
         enemy_vy_reg <= enemy_vy_next;
			
			enemyII_x_reg <= enemyII_x_next;
         enemyII_y_reg <= enemyII_y_next;
         enemyII_vx_reg <= enemyII_vx_next;
         enemyII_vy_reg <= enemyII_vy_next;
			
			enemyIII_x_reg <= enemyIII_x_next;
			enemyIII_y_reg <= enemyIII_y_next;
			enemyIII_vx_reg <= enemyIII_vx_next;
			enemyIII_vy_reg <= enemyIII_vy_next;
			
			shot_reg <= shot_next;
			rom_bit_player <= rom_next_player;
			btn_reg <= btn_next;
			arrow_reg <= arrow_next;
			
			rom_bit_enemy <= rom_next_enemy;
			rom_bit_enemyII <= rom_next_enemyII;
			rom_bit_enemyIII <= rom_next_enemyIII;
			contador <= contador_next;
			
      end if;
   end process;
	
	
	contador_next <=  std_logic_vector(unsigned(contador) + 1) when rst_enemy /= "110" else
							contador;
	
	-----------------------------------------------------------
	-- WALL
	-----------------------------------------------------------
   pix_x <= unsigned(pixel_x);
   pix_y <= unsigned(pixel_y);
   refr_tick <= '1' when (pix_y=481) and (pix_x=0) else
                '0';
   -- wall
   wall_on <=
      '1' when 	((zero<=pix_x) and (pix_x<=eight))
					or ((MAX_X-10<=pix_x) and (pix_x<=MAX_X))
					or ((zero<=pix_y) and (pix_y<=eight))
					or ((MAX_Y -33<=pix_y) and (pix_y<=MAX_Y))
					else
      '0';
   wall_rgb <= "001"; -- blue
	
	-----------------------------------------------------------
	-- CHESS
	-----------------------------------------------------------
	-- x -> 40,120,200,280,360,440,520,600
	-- y -> 30,90,150,210,270,330,390,450
--   chess_on <=
--      '1' when 	((1<=pix_x) and (pix_x<=39))
--					or ((121<=pix_x) and (pix_x<=159))
--					or ((201<=pix_x) and (pix_x<=239))
--					or ((281<=pix_x) and (pix_x<=319))
--					or ((361<=pix_x) and (pix_x<=399))
--					or ((441<=pix_x) and (pix_x<=479))
--					or ((521<=pix_x) and (pix_x<=559))
--					or ((601<=pix_x) and (pix_x<=639))
--					
--					or	((1<=pix_y) and (pix_y<=29))
--					or ((91<=pix_y) and (pix_y<=119))
--					or ((151<=pix_y) and (pix_y<=179))
--					or ((211<=pix_y) and (pix_y<=239))
--					or ((271<=pix_y) and (pix_y<=299))
--					or ((331<=pix_y) and (pix_y<=359))
--					or ((391<=pix_y) and (pix_y<=419))
--					--or ((450<=pix_y) and (pix_y<=479))
--					else
--      '0';
--   chess_rgb <= "000"; -- blue
	
	
	-----------------------------------------------------------	
	-- PLAYER
	-----------------------------------------------------------
	rom_addr_player <= pix_y(5 downto 0) - player_y_t(5 downto 0); --64 32 16 8 4 2 1
   rom_col_player <= pix_x(5 downto 0) - player_x_l(5 downto 0);
	
	--arrows 		btn
	--0 -> up		1
	--1 -> down		2
	--2 -> left		0
	--3 -> right	3
	--4 -> space
	
	process(btn, rom_bit_player, d_clr, btn_reg, arrows, arrow_reg)
   begin
		rom_next_player <= rom_bit_player;
		btn_next <= btn_reg;
		arrow_next <= arrow_reg;
      if d_clr='1'  then  --initial position of paddle
			rom_next_player <= PLAYER_ROM(to_integer(rom_addr_player), to_integer(rom_col_player));
      else
         if btn(2)='1' or arrows(1) = '1' then
				btn_next <= "0010";
				arrow_next <= "00010"; -- down 
				rom_next_player <= PLAYER_ROM(to_integer(rom_addr_player), to_integer(rom_col_player));
         elsif btn(1)='1' or arrows(0) = '1' then
				btn_next <= "0100";
				arrow_next <= "00001"; -- up
				rom_next_player <= PLAYER_ROM_BACK(to_integer(rom_addr_player), to_integer(rom_col_player));
			elsif btn(3)='1' or arrows(3) = '1'  then
				btn_next <= "1000";
				arrow_next <= "01000"; -- right
				rom_next_player <= PLAYER_ROM_SIDE(to_integer(rom_addr_player), to_integer(rom_col_player));
			elsif btn(0)='1' or arrows(2) = '1'  then
				btn_next <= "0001";
				arrow_next <= "00100"; -- left
				rom_next_player <= PLAYER_ROM_SIDE(to_integer(rom_addr_player), to_integer(not rom_col_player));	
			else
				--rom_next_player<= PLAYER_ROM(to_integer(rom_addr_player), to_integer(rom_col_player));--rom_next_player <= rom_bit_player;
				if btn_reg(1) ='1' or arrow_reg(0)='1' then -- up
					rom_next_player <= PLAYER_ROM(to_integer(rom_addr_player), to_integer(rom_col_player));
				elsif btn_reg(2) ='1' or arrow_reg(1)='1' then -- down
					rom_next_player <= PLAYER_ROM_BACK(to_integer(rom_addr_player), to_integer(rom_col_player));
				elsif btn_reg(3) ='1' or arrow_reg(3)='1' then -- right
					rom_next_player <= PLAYER_ROM_SIDE(to_integer(rom_addr_player), to_integer(rom_col_player));
				elsif btn_reg(0) = '1' or arrow_reg(2)='1' then -- left
					rom_next_player <= PLAYER_ROM_SIDE(to_integer(rom_addr_player), to_integer(not rom_col_player));
				end if;
				arrow_next <= "00000"; -- left
         end if;
      end if;
   end process;
	
	
   player_y_t <= player_y_reg;
	player_x_r <= player_x_reg;
   player_y_b <= player_y_t + ENEMY_SIZE - 1;
	player_x_l <= player_x_r + ENEMY_SIZE - 1;
   player_on <=
      '1' when (player_x_r<=pix_x) and (player_x_l>=pix_x) and
               (player_y_t<=pix_y) and (pix_y<=player_y_b) and (rom_bit_player/="000") else
      '0';
	player_rgb <= rom_bit_player;
	
   -- new player y and x-position
   process(btn,player_y_reg,player_y_b,player_y_t,refr_tick,gra_still,player_x_reg,player_x_r,
				player_x_l, d_clr, arrows, arrow_reg)
   begin
		player_y_next <= player_y_reg; -- no move
		player_x_next <= player_x_reg; -- no move
		
		if d_clr = '1' then  --initial position of paddle
			player_y_next <= to_unsigned((MAX_Y-ENEMY_SIZE)/2,10);
			player_x_next <= to_unsigned((MAX_X-ENEMY_SIZE)/2,10);
		elsif gra_still = '1' then 
			player_x_next <= player_x_reg;
			player_y_next <= player_y_reg;
		elsif refr_tick='1' then
			if (btn(2)='1' or arrow_reg(1)='1')and player_y_b<(MAX_Y-34-PLAYER_V) then --MAX_Y-33 -1-PLAYER_V
				player_y_next <= player_y_reg + PLAYER_V; -- move down
			elsif (btn(1)='1' or arrow_reg(0)='1')and player_y_t > (eight + PLAYER_V) then
				player_y_next <= player_y_reg - PLAYER_V; -- move up
			elsif (btn(3)='1' or arrow_reg(3)='1')and player_x_l <(MAX_X - 11 - PLAYER_V) then --MAX_X - 10 - PLAYER_V - 1
				player_x_next <= player_x_reg + PLAYER_V; -- move right
			elsif (btn(0)='1' or arrow_reg(2)='1')and player_x_r > (eight + PLAYER_V) then
				player_x_next <= player_x_reg - PLAYER_V; -- move left
			else 
				player_y_next <= player_y_reg; -- no move
				player_x_next <= player_x_reg; -- no move
			end if;
		end if;
   end process;
	
	-----------------------------------------------------------
	--BALL
	-----------------------------------------------------------
   -- square ball
   ball_x_l <= ball_x_reg; --ball_x_reg;
   ball_y_t <= ball_y_reg; --ball_y_reg;
   ball_x_r <= ball_x_l + 8 ;
   ball_y_b <= ball_y_t + 8 ;
--   sq_ball_on <=
--      '1' when (ball_x_l<=pix_x) and (pix_x<=ball_x_r) and
--               (ball_y_t<=pix_y) and (pix_y<=ball_y_b) else
--      '0';
   -- round ball
   rom_addr <= pix_y(2 downto 0) - ball_y_t(2 downto 0);
   rom_col <= pix_x(2 downto 0) - ball_x_l(2 downto 0);
   rom_data <= BALL_ROM(to_integer(rom_addr));
   rom_bit <= rom_data(to_integer(not rom_col));
   rd_ball_on <=
      '1' when (ball_x_l<=pix_x) and (pix_x<=ball_x_r) and
               (ball_y_t<=pix_y) and (pix_y<=ball_y_b) and 
					(rom_bit='1') 		and (player_on='0') else
      '0';
   ball_rgb <= "011";   -- cyan
   -- new ball position
   ball_x_next <=(player_x_reg + 16) when shot_reg = '0' else
		ball_x_reg + ball_vx_reg when refr_tick='1' else
      ball_x_reg;
   ball_y_next <=(player_y_reg + 16) when shot_reg = '0' else
		ball_y_reg + ball_vy_reg when refr_tick='1' else
      ball_y_reg;
   -- new ball velocity
   -- wuth new hit, miss signals
	
   process(ball_vx_reg,ball_vy_reg,ball_y_t,ball_x_l,ball_x_r,
           ball_y_t,ball_y_b,player_y_t,player_y_b,player_x_l, player_x_r,
			  rst_enemy, shot_reg, d_inc, shoot, btn_reg)
	begin
      --hit <='0';
      --miss <='0';
		shot_next <= shot_reg;
      ball_vx_next <= ball_vx_reg;
      ball_vy_next <= ball_vy_reg;
		if d_inc = '1' then		-- 00010 down 00001 up
			shot_next <= '0';
      elsif (shoot = '1' or arrows(4)='1') and (btn_reg(1) ='1' or arrow_reg(0)= '1') then            
			--UP
         ball_vx_next <= ENEMY_V_Z;
         ball_vy_next <= BALL_V_P;
			shot_next <= '1';
		elsif (shoot = '1' or arrows(4)='1')  and (btn_reg(2) ='1' or arrow_reg(1)= '1')  then          
         --DOWN
			ball_vx_next <= ENEMY_V_Z;
         ball_vy_next <= BALL_V_N;
			shot_next <= '1';
		elsif (shoot = '1' or arrows(4)='1')  and (btn_reg(3) ='1' or arrow_reg(3)= '1') then          
         --RIGHT
			ball_vx_next <= BALL_V_P;
         ball_vy_next <= ENEMY_V_Z;
			shot_next <= '1';
		elsif (shoot = '1' or arrows(4)='1')  and (btn_reg(0) ='1' or arrow_reg(2)= '1') then            
         --LEFT
			ball_vx_next <= BALL_V_N;
         ball_vy_next <= ENEMY_V_Z;
			shot_next <= '1';
      elsif ball_y_t < 1 or ball_y_b > (MAX_Y -33) or ball_x_l < 1 or (ball_x_r > (MAX_X -10)) then --paredes        		
			shot_next <= '0';
      end if;
   end process;
	
	
	-----------------------------------------------------------------------
	--ENEMY 
	-----------------------------------------------------------
	rom_addr_enemy <= pix_y(4 downto 1) - enemy_y_t(4 downto 1);
   rom_col_enemy <= pix_x(4 downto 1) - enemy_x_l(4 downto 1);
	
	-- enemy movement ------------
	process(enemy_vx_reg,enemy_vy_reg,enemy_y_t,enemy_x_l,enemy_x_r,
           enemy_y_b,player_y_t,player_y_b,gra_still,player_x_l, player_x_r, rom_next_enemy, rom_bit_enemy)
	begin
      enemy_vx_next <= enemy_vx_reg;
      enemy_vy_next <= enemy_vy_reg;
		rom_next_enemy <= rom_bit_enemy; 
		if gra_still='1' then            --initial velocity
         enemy_vx_next <= ENEMY_V_Z;
         enemy_vy_next <= ENEMY_V_Z;
			rom_next_enemy <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemy), to_integer(rom_col_enemy));
	
		elsif enemy_y_t = eight then  -- reach top border
         enemy_vy_next <= ENEMY_V_P;
			rom_next_enemy <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemy), to_integer(rom_col_enemy));
      elsif enemy_y_b = MAX_Y -33 then  -- reach bottom border
         enemy_vy_next <= enemy_V_N;
			rom_next_enemy <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemy), to_integer(rom_col_enemy));
      elsif enemy_x_l = eight  then -- reach left border
         enemy_vx_next <= enemy_V_P;
			rom_next_enemy <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemy), to_integer(rom_col_enemy));			
		elsif (enemy_x_r = MAX_X - 10) then-- reach right border
			enemy_vx_next <= enemy_V_N; 
			rom_next_enemy <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemy), to_integer(not rom_col_enemy));
		
		else
			if	enemy_y_t > player_y_b then -- bottom
				enemy_vy_next <= ENEMY_V_N;
			elsif enemy_y_b < player_y_t then-- top
				enemy_vy_next <= ENEMY_V_P;
			end if;
			if ( enemy_x_l >= (player_x_r - PLAYER_V) and enemy_x_r <= (player_x_l + PLAYER_V)) then --other
				enemy_vx_next <= ENEMY_V_Z;
				rom_next_enemy <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemy), to_integer(rom_col_enemy));
			elsif enemy_x_r < player_x_l then	-- left
				enemy_vx_next <= ENEMY_V_P;
				rom_next_enemy <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemy), to_integer(rom_col_enemy));
			elsif enemy_x_l > player_x_r then -- right
				enemy_vx_next <= ENEMY_V_N;
				rom_next_enemy <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemy), to_integer(not rom_col_enemy));
			end if;		
      end if;
   end process;
	
   enemy_x_l <= enemy_x_reg; --enemy_x_reg;
   enemy_y_t <= enemy_y_reg; --enemy_y_reg;
   enemy_x_r <= enemy_x_l + ENEMY_SIZE ;
   enemy_y_b <= enemy_y_t + ENEMY_SIZE ;
	enemy_on <=
      '1' when (enemy_x_l<=pix_x) and (enemy_x_r>=pix_x) and
               (enemy_y_t<=pix_y) and (pix_y<=enemy_y_b) and (rom_bit_enemy/="000") and 
					(rst_enemy = "010" or rst_enemy = "100" or rst_enemy = "110" or rst_enemy = "000")else
      '0';
	enemy_rgb <= rom_bit_enemy; 
	
   -- new enemy position--------------------
   enemy_x_next <=
		to_unsigned(eight,10) when gra_still='1' or 
						rst_enemy = "001" or rst_enemy = "011" or rst_enemy = "101" or rst_enemy = "111" else
		enemy_x_reg + enemy_vx_reg when refr_tick='1' else
      enemy_x_reg ;
		
   enemy_y_next <=
		to_unsigned(eight,10) when gra_still='1' or 
						rst_enemy = "001" or rst_enemy = "011" or rst_enemy = "101" or rst_enemy = "111" else
		enemy_y_reg + enemy_vy_reg when refr_tick='1' else
      enemy_y_reg ;
		
	--hiteI <= '0' when rst_enemy= "01";
	-----------------------------------------------------------------------
	--ENEMY 2
	-----------------------------------------------------------
	
	rom_addr_enemyII <= pix_y(4 downto 1) - enemyII_y_t(4 downto 1);
   rom_col_enemyII <= pix_x(4 downto 1) - enemyII_x_l(4 downto 1);
		
	-- enemyII movement ------------
	process(enemyII_vx_reg,enemyII_vy_reg,enemyII_y_t,enemyII_x_l,enemyII_x_r,
           enemyII_y_b,player_y_t,player_y_b,gra_still,player_x_l, player_x_r, rom_next_enemyII, rom_bit_enemyII)
	begin
      enemyII_vx_next <= enemyII_vx_reg;
      enemyII_vy_next <= enemyII_vy_reg;
		rom_next_enemyII <= rom_bit_enemyII; 
		if gra_still='1' then            --initial velocity
         enemyII_vx_next <= ENEMY_V_Z;
         enemyII_vy_next <= ENEMY_V_Z;
			rom_next_enemyII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyII), to_integer(not rom_col_enemyII));		
		elsif enemyII_y_t = eight then  -- reach top border
         enemyII_vy_next <= ENEMY_V_P;
			rom_next_enemyII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyII), to_integer(rom_col_enemyII));
      elsif enemyII_y_b = MAX_Y -33 then  -- reach bottom border
         enemyII_vy_next <= ENEMY_V_N;
			rom_next_enemyII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyII), to_integer(rom_col_enemyII));
      elsif enemyII_x_l = eight  then -- reach left border
         enemyII_vx_next <= ENEMY_V_N;
			rom_next_enemyII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyII), to_integer(rom_col_enemyII));			
		elsif (enemyII_x_r = MAX_X - 10) then-- reach right border
			enemyII_vx_next <= ENEMY_V_N; 
			rom_next_enemyII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyII), to_integer(not rom_col_enemyII));
			
		else
			if	enemyII_y_t > player_y_b then -- bottom
				enemyII_vy_next <= ENEMY_V_N;
			elsif enemyII_y_b < player_y_t then-- top
				enemyII_vy_next <= ENEMY_V_P;
			end if;
			if ( enemyII_x_l >= (player_x_r - PLAYER_V) and enemyII_x_r <= (player_x_l + PLAYER_V)) then --other
				enemyII_vx_next <= ENEMY_V_Z;
				rom_next_enemyII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyII), to_integer(rom_col_enemyII));
			elsif enemyII_x_r < player_x_l then	-- left
				enemyII_vx_next <= ENEMY_V_P;
				rom_next_enemyII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyII), to_integer(rom_col_enemyII));
			elsif enemyII_x_l > player_x_r then -- right
				enemyII_vx_next <= ENEMY_V_N;
				rom_next_enemyII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyII), to_integer(not rom_col_enemyII));
			else
				enemyII_vx_next <= ENEMY_V_N;
				enemyII_vy_next <= ENEMY_V_P;
				rom_next_enemyII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyII), to_integer(not rom_col_enemyII));
			end if;
      end if;
   end process;
	
	enemyII_x_l <= enemyII_x_reg; --ball_x_reg;
   enemyII_y_t <= enemyII_y_reg; --ball_y_reg;
   enemyII_x_r <= enemyII_x_l + ENEMY_SIZE ;
   enemyII_y_b <= enemyII_y_t + ENEMY_SIZE ;
	enemyII_on <=
      '1' when (enemyII_x_l<=pix_x) and (enemyII_x_r>=pix_x) and(enemyII_y_t<=pix_y) and (pix_y<=enemyII_y_b) and 
					(rom_bit_enemyII/="000") and (rst_enemy = "001" or rst_enemy = "100" or rst_enemy = "101" or rst_enemy = "000") else--and contador >= "01" else
      '0';
	enemyII_rgb <= rom_bit_enemyII; 
	
   -- new enemyII position--------------------
   enemyII_x_next <=
		to_unsigned((MAX_X -10 - ENEMY_SIZE),10) when gra_still='1' or 
						rst_enemy = "010" or rst_enemy = "011" or rst_enemy = "110" or rst_enemy = "111" else
		enemyII_x_reg + enemyII_vx_reg when refr_tick='1' else
      enemyII_x_reg ;
		
   enemyII_y_next <=
		to_unsigned(eight,10) when gra_still='1' or 
						rst_enemy = "010" or rst_enemy = "011" or rst_enemy = "110" or rst_enemy = "111" else
		enemyII_y_reg + enemyII_vy_reg when refr_tick='1' else
      enemyII_y_reg ;

	--hiteII <= '0' when rst_enemy= "10";
	-----------------------------------------------------------------------
	--ENEMY 3
	-----------------------------------------------------------

	rom_addr_enemyIII <= pix_y(4 downto 1) - enemyIII_y_t(4 downto 1);
   rom_col_enemyIII <= pix_x(4 downto 1) - enemyIII_x_l(4 downto 1);
		
	-- enemyIII movement ------------
	process(enemyIII_vx_reg,enemyIII_vy_reg,enemyIII_y_t,enemyIII_x_l,enemyIII_x_r,
           enemyIII_y_b,player_y_t,player_y_b,gra_still,player_x_l, player_x_r, rom_next_enemyIII, rom_bit_enemyIII)
	begin
      enemyIII_vx_next <= enemyIII_vx_reg;
      enemyIII_vy_next <= enemyIII_vy_reg;
		rom_next_enemyIII <= rom_bit_enemyIII; 
		if gra_still='1' then            --initial velocity
         enemyIII_vx_next <= ENEMY_V_Z;
         enemyIII_vy_next <= ENEMY_V_Z;
			rom_next_enemyIII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyIII), to_integer(not rom_col_enemyIII));			
		elsif enemyIII_y_t = eight then  -- reach top border
         enemyIII_vy_next <= ENEMY_V_P;
			rom_next_enemyIII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyIII), to_integer(rom_col_enemyIII));
      elsif enemyIII_y_b = MAX_Y -33 then  -- reach bottom border
         enemyIII_vy_next <= ENEMY_V_N;
			rom_next_enemyIII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyIII), to_integer(rom_col_enemyIII));
      elsif enemyIII_x_l = eight  then -- reach left border
         enemyIII_vx_next <= ENEMY_V_N;
			rom_next_enemyIII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyIII), to_integer(rom_col_enemyIII));			
		elsif (enemyIII_x_r = MAX_X -10) then-- reach right border
			enemyIII_vx_next <= ENEMY_V_N; 
			rom_next_enemyIII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyIII), to_integer(not rom_col_enemyIII));
			
		else
			if	enemyIII_y_t > player_y_b then -- bottom
				enemyIII_vy_next <= ENEMY_V_N;
			elsif enemyIII_y_b < player_y_t then-- top
				enemyIII_vy_next <= ENEMY_V_P;
			end if;
			if ( enemyIII_x_l >= (player_x_r - PLAYER_V) and enemyIII_x_r <= (player_x_l + PLAYER_V)) then --other
				enemyIII_vx_next <= ENEMY_V_Z;
				rom_next_enemyIII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyIII), to_integer(rom_col_enemyIII));
			elsif enemyIII_x_r < player_x_l then	-- left
				enemyIII_vx_next <= ENEMY_V_P;
				rom_next_enemyIII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyIII), to_integer(rom_col_enemyIII));
			elsif enemyIII_x_l > player_x_r then -- right
				enemyIII_vx_next <= ENEMY_V_N;
				rom_next_enemyIII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyIII), to_integer(not rom_col_enemyIII));
			else
				enemyIII_vx_next <= ENEMY_V_N;
				enemyIII_vy_next <= ENEMY_V_N;
				rom_next_enemyIII <= ENEMY_ROM_SIDE(to_integer(rom_addr_enemyIII), to_integer(not rom_col_enemyIII));
			end if;
      end if;
   end process;
	
	enemyIII_x_l <= enemyIII_x_reg; --ball_x_reg;
   enemyIII_y_t <= enemyIII_y_reg; --ball_y_reg;
   enemyIII_x_r <= enemyIII_x_l + ENEMY_SIZE ;
   enemyIII_y_b <= enemyIII_y_t + ENEMY_SIZE ;
	enemyIII_on <=
      '1' when (enemyIII_x_l<=pix_x) and (enemyIII_x_r>=pix_x) and(enemyIII_y_t<=pix_y) and (pix_y<=enemyIII_y_b) and 
					(rom_bit_enemyIII/="000") and (rst_enemy = "000" or rst_enemy = "001" or rst_enemy = "010" or rst_enemy = "011") else--and contador >= "01" else
      '0';
	enemyIII_rgb <= rom_bit_enemyIII; 
	
   -- new enemyIII position--------------------
   enemyIII_x_next <=
		to_unsigned((MAX_X/2),10) when gra_still='1' or 
						rst_enemy = "100" or rst_enemy = "101" or rst_enemy = "110" or rst_enemy = "111" else
		enemyIII_x_reg + enemyIII_vx_reg when refr_tick='1' else
      enemyIII_x_reg ;
		
   enemyIII_y_next <=
		to_unsigned((MAX_Y -33 - ENEMY_SIZE),10) when gra_still='1' or
						rst_enemy = "100" or rst_enemy = "101" or rst_enemy = "110" or rst_enemy = "111" else
		enemyIII_y_reg + enemyIII_vy_reg when refr_tick='1' else
      enemyIII_y_reg ;

	---hiteIII <= '0' when rst_enemy= "11";
	
	-----------------------------------------------------------
	
--	process(enemy_on, enemyII_on, enemyIII_on, rd_ball_on, player_on, rst_enemy)
--	begin
--		
--		hiteI <='0';
--		hiteII <= '0';
--		hiteIII <= '0';
--		
--		if rst_enemy(0) = '1' then
--			hiteI <= '0';
--		elsif rst_enemy(1) = '1' then
--			hiteII <= '0';
--		elsif rst_enemy(2) = '1' then
--			hiteIII <= '0';
--		end if;
--	end process;
	-----------------------------------------------------------	
   -- rgb multiplexing circuit
	-----------------------------------------------------------
   process(	wall_on,rd_ball_on,wall_rgb,player_rgb,ball_rgb,
				enemy_on, enemy_rgb, enemyII_on, enemyII_rgb,
				player_on, enemyIII_on, enemyIII_rgb)
   begin
		miss <= '0';
		hiteI <= '0';
		hiteII <= '0';
		hiteIII <= '0';
			
		if (player_on = '1') and ((enemy_on = '1') or (enemyII_on = '1') or (enemyIII_on = '1')) then
			miss <='1';
		elsif (rd_ball_on = '1') and (enemy_on = '1') then
			hiteI <= '1';
		elsif (rd_ball_on = '1') and (enemyII_on = '1') then
			hiteII <= '1';
		elsif (rd_ball_on = '1') and (enemyIII_on = '1') then
			hiteIII <= '1';
			
      elsif wall_on='1' then
         rgb <= wall_rgb;
      elsif player_on='1' then
         rgb <= player_rgb;
		elsif enemy_on ='1' then 
			rgb <= enemy_rgb;
		elsif enemyII_on ='1' then 
			rgb <= enemyII_rgb;
		elsif enemyIII_on ='1' then 
			rgb <= enemyIII_rgb;
      elsif rd_ball_on='1' then
         rgb <= ball_rgb;
--		elsif chess_on='1' then
--         rgb <= chess_rgb;
			--rgb <= "101";
      else
			hiteI <= '0';
			hiteII <= '0';
			hiteIII <= '0';
         rgb <= "111"; -- yellow background
      end if;
   end process;
   -- new graphic_on signal
   graph_on <= wall_on or player_on or rd_ball_on or enemy_on or enemyII_on or enemyIII_on;
end arch;
